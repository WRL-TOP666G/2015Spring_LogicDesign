module adder_32bit(in1, in2, sum);
	input [31:0]in1, in2;
	output [31:0]sum;
	
	/* design here */
	
endmodule
