module ALU_3(A,B,S,C_2,F,G,P,C_3);
  input  [11:8]A;
  input  [11:8]B;
  input  [2:0]S;
  input  C_2;
  output signed [11:8]F;
  output G,P,C_3;
  reg signed   [11:8]F;
  reg    C_3;
  reg    G,P;
  
  always@(C_2,G,P) 
   begin
    C_3=G+P*C_2;
   
   end
 always@(S or A or B)
 begin
   case(S)
     3'b000: begin F=4'b0000  ;G=1'b1       ;P=1'b1    ; end
     3'b001: begin F=B-A      ;G=~(~A&~B|A) ;P=~(A&~B) ; end
     3'b010: begin F=A-B      ;G=~(~A|A&B)  ;P=~(~A&B) ; end
     3'b011: begin F=A+B      ;G=~(~A|A&~B) ;P=~(~A&~B); end
     3'b100: begin F=A^B      ;G=~(A^B)     ;P=~(~A&B) ; end
     3'b101: begin F=A|B      ;G=~(A|B)     ;P=~(A^B)  ; end
     3'b110: begin F=A&B      ;G=~B         ;P=~(~A&B) ; end
     3'b111: begin F=4'b1111  ;G=1'b0       ;P=(A&B)   ; end
   endcase
 end
 
 

  
   
   
endmodule
