module program_counter(clk, rst, next_pc, pc);
	input clk, rst;
	input [31:0]next_pc;
	output [31:0]pc;
	
	/* design here */
	
endmodule
